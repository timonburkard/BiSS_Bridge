library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_data_checker is
end tb_data_checker;

architecture tb of tb_data_checker is
    -- Generics and constants
    constant CLK_PERIOD : time := 8 ns;  -- 125 MHz
    constant DATA_WIDTH : integer := 22;
    constant CRC_WIDTH  : integer := 6;

    -- Signals
    signal clk           : STD_LOGIC := '0';
    signal rst           : STD_LOGIC := '1';
    signal position_raw  : STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0) := (others => '0');
    signal crc           : STD_LOGIC_VECTOR(CRC_WIDTH-1 downto 0) := (others => '0');
    signal position      : STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
    signal error_bit     : STD_LOGIC := '0';
    signal warning_bit   : STD_LOGIC := '0';
    signal crc_fail_bit  : STD_LOGIC;
    signal data_valid_out : STD_LOGIC;

    -- Hard-coded test vectors with pre-calculated CRC values (now includes status bits)
    type test_vector_t is record
        position : STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
        crc      : STD_LOGIC_VECTOR(CRC_WIDTH-1 downto 0);
        error    : STD_LOGIC;  -- decoded error (active-high)
        warning  : STD_LOGIC;  -- decoded warning (active-high)
    end record;

    type test_vector_array_t is array (natural range <>) of test_vector_t;

    -- Test vectors generated by 6_tools/calculate_crc.py (includes E/W bits in CRC)
    constant TEST_VECTORS : test_vector_array_t := (
        (position => "0000000000000000000000", crc => "111010", error => '0', warning => '0'),  -- All zeros
        (position => "1111111111111111111111", crc => "101111", error => '0', warning => '0'),  -- All ones (22-bit)
        (position => "0100100011010001010110", crc => "110101", error => '0', warning => '0'),  -- Test pattern 1
        (position => "1010111100110111101111", crc => "010000", error => '0', warning => '0'),  -- Test pattern 2
        (position => "0101010100001100100001", crc => "110110", error => '0', warning => '0'),  -- Test pattern 3
        (position => "1111101101110010111010", crc => "011000", error => '0', warning => '0'),  -- Test pattern 4
        (position => "0000101110111111001010", crc => "011100", error => '0', warning => '0'),  -- Test pattern real
        (position => "0000010010001101000101", crc => "001011", error => '1', warning => '0'),  -- Error=1, Warning=0
        (position => "0000010010001101000101", crc => "001110", error => '0', warning => '1')   -- Error=0, Warning=1
    );

begin

    -- Instantiate DUT
    DUT : entity work.Data_Checker
        generic map (
            DATA_WIDTH => DATA_WIDTH,
            CRC_WIDTH  => CRC_WIDTH
        )
        port map (
            clk          => clk,
            rst          => rst,
            position_raw => position_raw,
            crc          => crc,
            error_bit    => error_bit,
            warning_bit  => warning_bit,
            data_valid_in => '1',
            position     => position,
            data_valid_out => data_valid_out,
            crc_fail_bit => crc_fail_bit
        );

    -- Clock generation
    clk_process : process
    begin
        wait for CLK_PERIOD / 2;
        clk <= not clk;
    end process;

    -- Main test process
    test_process : process
        variable test_idx : integer;
    begin
        -- Reset
        rst <= '1';
        wait for 5 * CLK_PERIOD;
        rst <= '0';
        wait for CLK_PERIOD;

        -- Test 1: Valid data with correct CRC from test vectors
        report "TEST 1: Valid position data with correct CRC";
        position_raw <= TEST_VECTORS(2).position;
        crc <= TEST_VECTORS(2).crc;
        error_bit   <= TEST_VECTORS(2).error;
        warning_bit <= TEST_VECTORS(2).warning;

        wait for 2 * CLK_PERIOD;

        assert position = TEST_VECTORS(2).position
            report "ERROR: Position should be latched"
            severity ERROR;
        assert crc_fail_bit = '0'
            report "ERROR: CRC should be valid (crc_fail_bit should be 0)"
            severity ERROR;

        report "TEST 1: PASSED - Valid data accepted";

        -- Test 2: Invalid CRC
        report "TEST 2: Invalid CRC detection";
        position_raw <= TEST_VECTORS(3).position;
        crc <= "000000";  -- Wrong CRC
        error_bit   <= TEST_VECTORS(3).error;
        warning_bit <= TEST_VECTORS(3).warning;

        wait for 2 * CLK_PERIOD;

        assert crc_fail_bit = '1'
            report "ERROR: CRC should be invalid (crc_fail_bit should be 1)"
            severity ERROR;

        report "TEST 2: PASSED - Invalid CRC detected";

        -- Test 3: Error bit coverage
        report "TEST 3: Error bit in CRC coverage";
        position_raw <= TEST_VECTORS(7).position;  -- Same position, error=1
        crc <= TEST_VECTORS(7).crc;  -- Different CRC due to error bit
        error_bit   <= TEST_VECTORS(7).error;
        warning_bit <= TEST_VECTORS(7).warning;

        wait for 2 * CLK_PERIOD;

        assert crc_fail_bit = '0'
            report "ERROR: CRC with error=1 should be valid"
            severity ERROR;

        report "TEST 3: PASSED - Error bit correctly included in CRC";

        -- Test 4: Warning bit coverage
        report "TEST 4: Warning bit in CRC coverage";
        position_raw <= TEST_VECTORS(8).position;  -- Same position, warning=1
        crc <= TEST_VECTORS(8).crc;  -- Different CRC due to warning bit
        error_bit   <= TEST_VECTORS(8).error;
        warning_bit <= TEST_VECTORS(8).warning;

        wait for 2 * CLK_PERIOD;

        assert crc_fail_bit = '0'
            report "ERROR: CRC with warning=1 should be valid"
            severity ERROR;

        report "TEST 4: PASSED - Warning bit correctly included in CRC";

        -- Test 5: All test vectors
        report "TEST 5: Testing all predefined test vectors";
        for i in TEST_VECTORS'range loop
            position_raw <= TEST_VECTORS(i).position;
            crc <= TEST_VECTORS(i).crc;
            error_bit   <= TEST_VECTORS(i).error;
            warning_bit <= TEST_VECTORS(i).warning;

            wait for 2 * CLK_PERIOD;

            assert position = TEST_VECTORS(i).position
                report "ERROR: Position mismatch at vector " & integer'image(i)
                severity ERROR;
            assert crc_fail_bit = '0'
                report "ERROR: CRC should be valid for vector " & integer'image(i)
                severity ERROR;

            report "  Vector " & integer'image(i) & ": position = " &
                   integer'image(TO_INTEGER(UNSIGNED(position))) &
                   ", crc = " & integer'image(TO_INTEGER(UNSIGNED(TEST_VECTORS(i).crc))) &
                   ", E=" & STD_LOGIC'image(TEST_VECTORS(i).error) &
                   ", W=" & STD_LOGIC'image(TEST_VECTORS(i).warning) & " - OK";
        end loop;

        report "TEST 5: PASSED - All test vectors passed CRC validation";

        -- Test complete
        report "All tests completed successfully";
        wait;

    end process;

end tb;
