library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package biss_bridge_pkg is
  constant C_CLK_FREQ_HZ : positive := 125_000_000; -- clock frequency
end;
